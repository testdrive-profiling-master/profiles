module TOP # ( 
	parameter	DATA_WIDTH
) (
	input		CLK,
	input		nRE,
	input		nCLR,
	input		nWE,
	input [31:0]		DIN,
	output [31:0]		DOUT
);

endmodule
