`include "DUTs/processor_axi_wrapper/includes.vh"
`include "DUTs/processor_axi_wrapper/processor_top.v"

module dut_wrapper_v1_0 #(
	parameter			C_CLKIN_PERIOD			= 4,
	// AXI_LITE
	parameter integer	C_M_AXILITE_ADDR_WIDTH	= 20,
	// M_AXI
	parameter integer	C_M_AXI_ID_WIDTH		= 1,
	parameter integer	C_M_AXI_ADDR_WIDTH		= 32,
	parameter integer	C_M_AXI_DATA_WIDTH		= 512
) (
	//// system
	input									ACLK,
	input									nRST,
	output									INTR,

	//// slave APB -------------------------
	input									S_PSEL,
	input									S_PENABLE,
	input									S_PWRITE,
	input	[15:0]							S_PADDR,
	input	[31:0]							S_PWDATA,
	output	[31:0]							S_PRDATA,
	output									S_PREADY,
	output									S_PSLVERR,

	//// external control AXI_LITE ---------
	// write address
	output	[C_M_AXILITE_ADDR_WIDTH-1 : 0]	EX_AWADDR,
	output									EX_AWVALID,
	input									EX_AWREADY,
	// write data
	output	[31 : 0]						EX_WDATA,
	output	[3 : 0]							EX_WSTRB,
	output									EX_WVALID,
	input									EX_WREADY,
	// read address
	output	[C_M_AXILITE_ADDR_WIDTH-1 : 0]	EX_ARADDR,
	output									EX_ARVALID,
	input									EX_ARREADY,
	// read data
	input	[31 : 0]						EX_RDATA,
	input	[1 : 0]							EX_RRESP,
	input									EX_RVALID,
	output									EX_RREADY,
	// bus
	input	[1 : 0]							EX_BRESP,
	input									EX_BVALID,
	output									EX_BREADY,

	//// master AXI_0 ----------------------
	// write address
	output	[C_M_AXI_ID_WIDTH-1 : 0]		M0_AWID,
	output	[C_M_AXI_ADDR_WIDTH-1 : 0]		M0_AWADDR,
	output	[7 : 0]							M0_AWLEN,
	output	[2 : 0]							M0_AWSIZE,
	output	[1 : 0]							M0_AWBURST,
	output									M0_AWLOCK,
	output	[3 : 0]							M0_AWCACHE,
	output	[2 : 0]							M0_AWPROT,
	output	[3 : 0]							M0_AWREGION,
	output	[3 : 0]							M0_AWQOS,
	output									M0_AWVALID,
	input									M0_AWREADY,
	// write data
	output	[C_M_AXI_ID_WIDTH-1 : 0]		M0_WID,
	output	[C_M_AXI_DATA_WIDTH-1 : 0]		M0_WDATA,
	output	[C_M_AXI_DATA_WIDTH/8-1 : 0]	M0_WSTRB,
	output									M0_WLAST,
	output									M0_WVALID,
	input									M0_WREADY,
	// read address
	output	[C_M_AXI_ID_WIDTH-1 : 0]		M0_ARID,
	output	[C_M_AXI_ADDR_WIDTH-1 : 0]		M0_ARADDR,
	output	[7 : 0]							M0_ARLEN,
	output	[2 : 0]							M0_ARSIZE,
	output	[1 : 0]							M0_ARBURST,
	output									M0_ARLOCK,
	output	[3 : 0]							M0_ARCACHE,
	output	[2 : 0]							M0_ARPROT,
	output	[3 : 0]							M0_ARREGION,
	output	[3 : 0]							M0_ARQOS,
	output									M0_ARVALID,
	input									M0_ARREADY,
	// read data
	input	[C_M_AXI_ID_WIDTH-1 : 0]		M0_RID,
	input	[C_M_AXI_DATA_WIDTH-1 : 0]		M0_RDATA,
	input	[1 : 0]							M0_RRESP,
	input									M0_RLAST,
	input									M0_RVALID,
	output									M0_RREADY,
	// bus
	input	[C_M_AXI_ID_WIDTH-1 : 0]		M0_BID,
	input	[1 : 0]							M0_BRESP,
	input									M0_BVALID,
	output									M0_BREADY,
	
	//// master AXI_0 ----------------------
	// write address
	output	[C_M_AXI_ID_WIDTH-1 : 0]		M1_AWID,
	output	[C_M_AXI_ADDR_WIDTH-1 : 0]		M1_AWADDR,
	output	[7 : 0]							M1_AWLEN,
	output	[2 : 0]							M1_AWSIZE,
	output	[1 : 0]							M1_AWBURST,
	output									M1_AWLOCK,
	output	[3 : 0]							M1_AWCACHE,
	output	[2 : 0]							M1_AWPROT,
	output	[3 : 0]							M1_AWREGION,
	output	[3 : 0]							M1_AWQOS,
	output									M1_AWVALID,
	input									M1_AWREADY,
	// write data
	output	[C_M_AXI_ID_WIDTH-1 : 0]		M1_WID,
	output	[C_M_AXI_DATA_WIDTH-1 : 0]		M1_WDATA,
	output	[C_M_AXI_DATA_WIDTH/8-1 : 0]	M1_WSTRB,
	output									M1_WLAST,
	output									M1_WVALID,
	input									M1_WREADY,
	// read address
	output	[C_M_AXI_ID_WIDTH-1 : 0]		M1_ARID,
	output	[C_M_AXI_ADDR_WIDTH-1 : 0]		M1_ARADDR,
	output	[7 : 0]							M1_ARLEN,
	output	[2 : 0]							M1_ARSIZE,
	output	[1 : 0]							M1_ARBURST,
	output									M1_ARLOCK,
	output	[3 : 0]							M1_ARCACHE,
	output	[2 : 0]							M1_ARPROT,
	output	[3 : 0]							M1_ARREGION,
	output	[3 : 0]							M1_ARQOS,
	output									M1_ARVALID,
	input									M1_ARREADY,
	// read data
	input	[C_M_AXI_ID_WIDTH-1 : 0]		M1_RID,
	input	[C_M_AXI_DATA_WIDTH-1 : 0]		M1_RDATA,
	input	[1 : 0]							M1_RRESP,
	input									M1_RLAST,
	input									M1_RVALID,
	output									M1_RREADY,
	// bus
	input	[C_M_AXI_ID_WIDTH-1 : 0]		M1_BID,
	input	[1 : 0]							M1_BRESP,
	input									M1_BVALID,
	output									M1_BREADY
);

// implementation ------------------------------------------------------------
// DUT processor
processor_axi_wrapper #(
	.C_CLKIN_PERIOD			(C_CLKIN_PERIOD),
	.C_M_AXILITE_ADDR_WIDTH	(C_M_AXILITE_ADDR_WIDTH),
	.C_M_AXI_ID_WIDTH		(C_M_AXI_ID_WIDTH),
	.C_M_AXI_ADDR_WIDTH		(C_M_AXI_ADDR_WIDTH),
	.C_M_AXI_DATA_WIDTH		(C_M_AXI_DATA_WIDTH)
) processor_inst (
	//// system
	.CLK			(ACLK),
	.nRST			(nRST),
	.INTR			(INTR),
	//// slave APB -------------------------
	.S_PSEL			(S_PSEL),
	.S_PENABLE		(S_PENABLE),
	.S_PWRITE		(S_PWRITE),
	.S_PADDR		(S_PADDR),
	.S_PWDATA		(S_PWDATA),
	.S_PRDATA		(S_PRDATA),
	.S_PREADY		(S_PREADY),
	.S_PSLVERR		(S_PSLVERR),
	//// external control AXI_LITE ---------
	.EX_AWADDR		(EX_AWADDR),
	.EX_AWVALID		(EX_AWVALID),
	.EX_AWREADY		(EX_AWREADY),
	.EX_WDATA		(EX_WDATA),
	.EX_WSTRB		(EX_WSTRB),
	.EX_WVALID		(EX_WVALID),
	.EX_WREADY		(EX_WREADY),
	.EX_ARADDR		(EX_ARADDR),
	.EX_ARVALID		(EX_ARVALID),
	.EX_ARREADY		(EX_ARREADY),
	.EX_RDATA		(EX_RDATA),
	.EX_RRESP		(EX_RRESP),
	.EX_RVALID		(EX_RVALID),
	.EX_RREADY		(EX_RREADY),
	.EX_BRESP		(EX_BRESP),
	.EX_BVALID		(EX_BVALID),
	.EX_BREADY		(EX_BREADY),
	//// AXI master #0 interface ------------
	.M0_AWID		(M0_AWID),
	.M0_AWADDR		(M0_AWADDR),
	.M0_AWLEN		(M0_AWLEN),
	.M0_AWSIZE		(M0_AWSIZE),
	.M0_AWBURST		(M0_AWBURST),
	.M0_AWLOCK		(M0_AWLOCK),
	.M0_AWCACHE		(M0_AWCACHE),
	.M0_AWPROT		(M0_AWPROT),
	.M0_AWREGION	(M0_AWREGION),
	.M0_AWQOS		(M0_AWQOS),
	.M0_AWVALID		(M0_AWVALID),
	.M0_AWREADY		(M0_AWREADY),
	.M0_WID			(M0_WID),
	.M0_WDATA		(M0_WDATA),
	.M0_WSTRB		(M0_WSTRB),
	.M0_WLAST		(M0_WLAST),
	.M0_WVALID		(M0_WVALID),
	.M0_WREADY		(M0_WREADY),
	.M0_BID			(M0_BID),
	.M0_BRESP		(M0_BRESP),
	.M0_BVALID		(M0_BVALID),
	.M0_BREADY		(M0_BREADY),
	.M0_ARID		(M0_ARID),
	.M0_ARADDR		(M0_ARADDR),
	.M0_ARLEN		(M0_ARLEN),
	.M0_ARSIZE		(M0_ARSIZE),
	.M0_ARBURST		(M0_ARBURST),
	.M0_ARLOCK		(M0_ARLOCK),
	.M0_ARCACHE		(M0_ARCACHE),
	.M0_ARPROT		(M0_ARPROT),
	.M0_ARREGION	(M0_ARREGION),
	.M0_ARQOS		(M0_ARQOS),
	.M0_ARVALID		(M0_ARVALID),
	.M0_ARREADY		(M0_ARREADY),
	.M0_RID			(M0_RID),
	.M0_RDATA		(M0_RDATA),
	.M0_RRESP		(M0_RRESP),
	.M0_RLAST		(M0_RLAST),
	.M0_RVALID		(M0_RVALID),
	.M0_RREADY		(M0_RREADY),
	//// AXI master #1 interface ------------
	.M1_AWID		(M1_AWID),
	.M1_AWADDR		(M1_AWADDR),
	.M1_AWLEN		(M1_AWLEN),
	.M1_AWSIZE		(M1_AWSIZE),
	.M1_AWBURST		(M1_AWBURST),
	.M1_AWLOCK		(M1_AWLOCK),
	.M1_AWCACHE		(M1_AWCACHE),
	.M1_AWPROT		(M1_AWPROT),
	.M1_AWREGION	(M1_AWREGION),
	.M1_AWQOS		(M1_AWQOS),
	.M1_AWVALID		(M1_AWVALID),
	.M1_AWREADY		(M1_AWREADY),
	.M1_WID			(M1_WID),
	.M1_WDATA		(M1_WDATA),
	.M1_WSTRB		(M1_WSTRB),
	.M1_WLAST		(M1_WLAST),
	.M1_WVALID		(M1_WVALID),
	.M1_WREADY		(M1_WREADY),
	.M1_BID			(M1_BID),
	.M1_BRESP		(M1_BRESP),
	.M1_BVALID		(M1_BVALID),
	.M1_BREADY		(M1_BREADY),
	.M1_ARID		(M1_ARID),
	.M1_ARADDR		(M1_ARADDR),
	.M1_ARLEN		(M1_ARLEN),
	.M1_ARSIZE		(M1_ARSIZE),
	.M1_ARBURST		(M1_ARBURST),
	.M1_ARLOCK		(M1_ARLOCK),
	.M1_ARCACHE		(M1_ARCACHE),
	.M1_ARPROT		(M1_ARPROT),
	.M1_ARREGION	(M1_ARREGION),
	.M1_ARQOS		(M1_ARQOS),
	.M1_ARVALID		(M1_ARVALID),
	.M1_ARREADY		(M1_ARREADY),
	.M1_RID			(M1_RID),
	.M1_RDATA		(M1_RDATA),
	.M1_RRESP		(M1_RRESP),
	.M1_RLAST		(M1_RLAST),
	.M1_RVALID		(M1_RVALID),
	.M1_RREADY		(M1_RREADY)
);

endmodule
