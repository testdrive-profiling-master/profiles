//================================================================================
// Copyright (c) 2013 ~ 2019. HyungKi Jeong(clonextop@gmail.com)
// All rights reserved.
// 
// The 3-Clause BSD License (https://opensource.org/licenses/BSD-3-Clause)
// 
// Redistribution and use in source and binary forms,
// with or without modification, are permitted provided
// that the following conditions are met:
// 
// 1. Redistributions of source code must retain the above copyright notice,
//    this list of conditions and the following disclaimer.
// 
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
// 
// 3. Neither the name of the copyright holder nor the names of its contributors
//    may be used to endorse or promote products derived from this software
//    without specific prior written permission.
// 
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
// THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
// PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS
// BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE
// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
// HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
// STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN
// ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY
// OF SUCH DAMAGE.
// 
// Title : Meitner processor v1.1
// Rev.  : 10/31/2019 Thu (clonextop@gmail.com)
//================================================================================
`include "MTSP_Defines.vh"

module MTSP_SF_RSQ_LUT(CLK, index, REF);
// port definition -----------------------------------------------------------
input	CLK;
input	[7:0]		index;		// LUT index
output reg	[31:0]	REF;		// Reference Value

// register definition & assignment ------------------------------------------

// behavior code -------------------------------------------------------------
`ALWAYS_CLOCK begin
	case(index) //		 Reference Reference^3/2						 x.xxx...   0.0xxx...             x.xxx...   0.0xxx...
		0 :
			REF <= 32'b1000011110000000_1011001111110110;	//									Odd   0 : 1.0585946, 0.3514919
		1 :
			REF <= 32'b1011111110100000_1111111010000001;	//Even   0 : 1.4970789, 0.4970846
		2 :
			REF <= 32'b1000011011111001_1011000111100010;	//									Odd   1 : 1.0544995, 0.3474284
		3 :
			REF <= 32'b1011111011100010_1111101110010000;	//Even   1 : 1.4912875, 0.4913380
		4 :
			REF <= 32'b1000011001110101_1010111111010111;	//									Odd   2 : 1.0504515, 0.3434426
		5 :
			REF <= 32'b1011111000100110_1111100010101101;	//Even   2 : 1.4855627, 0.4857012
		6 :
			REF <= 32'b1000010111110010_1010110111010111;	//									Odd   3 : 1.0464498, 0.3395325
		7 :
			REF <= 32'b1011110101101101_1111010111011001;	//Even   3 : 1.4799033, 0.4801714
		8 :
			REF <= 32'b1000010101110000_1010101111100000;	//									Odd   4 : 1.0424933, 0.3356960
		9 :
			REF <= 32'b1011110010110110_1111001100010001;	//Even   4 : 1.4743083, 0.4747458
		10 :
			REF <= 32'b1000010011110000_1010100111110010;	//									Odd   5 : 1.0385816, 0.3319312
		11 :
			REF <= 32'b1011110000000000_1111000001011000;	//Even   5 : 1.4687761, 0.4694216
		12 :
			REF <= 32'b1000010001110001_1010100000001110;	//									Odd   6 : 1.0347135, 0.3282363
		13 :
			REF <= 32'b1011101101001101_1110110110101011;	//Even   6 : 1.4633058, 0.4641961
		14 :
			REF <= 32'b1000001111110100_1010011000110011;	//									Odd   7 : 1.0308883, 0.3246093
		15 :
			REF <= 32'b1011101010011100_1110101100001010;	//Even   7 : 1.4578962, 0.4590669
		16 :
			REF <= 32'b1000001101111000_1010010001100000;	//									Odd   8 : 1.0271052, 0.3210487
		17 :
			REF <= 32'b1011100111101101_1110100001110110;	//Even   8 : 1.4525461, 0.4540315
		18 :
			REF <= 32'b1000001011111101_1010001010010110;	//									Odd   9 : 1.0233635, 0.3175528
		19 :
			REF <= 32'b1011100100111111_1110010111101110;	//Even   9 : 1.4472544, 0.4490874
		20 :
			REF <= 32'b1000001010000100_1010000011010100;	//									Odd  10 : 1.0196623, 0.3141198
		21 :
			REF <= 32'b1011100010010100_1110001101110010;	//Even  10 : 1.4420203, 0.4442325
		22 :
			REF <= 32'b1000001000001100_1001111100011010;	//									Odd  11 : 1.0160010, 0.3107482
		23 :
			REF <= 32'b1011011111101010_1110000100000001;	//Even  11 : 1.4368424, 0.4394644
		24 :
			REF <= 32'b1000000110010101_1001110101101000;	//									Odd  12 : 1.0123789, 0.3074365
		25 :
			REF <= 32'b1011011101000010_1101111010011011;	//Even  12 : 1.4317200, 0.4347809
		26 :
			REF <= 32'b1000000100100000_1001101110111101;	//									Odd  13 : 1.0087953, 0.3041832
		27 :
			REF <= 32'b1011011010011100_1101110001000000;	//Even  13 : 1.4266520, 0.4301801
		28 :
			REF <= 32'b1000000010101100_1001101000011010;	//									Odd  14 : 1.0052494, 0.3009869
		29 :
			REF <= 32'b1011010111111000_1101100111110000;	//Even  14 : 1.4216373, 0.4256598
		30 :
			REF <= 32'b1000000000111001_1001100001111111;	//									Odd  15 : 1.0017407, 0.2978462
		31 :
			REF <= 32'b1011010101010101_1101011110101001;	//Even  15 : 1.4166752, 0.4212182
		32 :
			REF <= 32'b0111111111000111_1001011011101010;	//									Odd  16 : 0.9982684, 0.2947598
		33 :
			REF <= 32'b1011010010110100_1101010101101101;	//Even  16 : 1.4117647, 0.4168532
		34 :
			REF <= 32'b0111111101010110_1001010101011101;	//									Odd  17 : 0.9948320, 0.2917262
		35 :
			REF <= 32'b1011010000010101_1101001100111011;	//Even  17 : 1.4069049, 0.4125632
		36 :
			REF <= 32'b0111111011100111_1001001111010110;	//									Odd  18 : 0.9914309, 0.2887444
		37 :
			REF <= 32'b1011001101110111_1101000100010010;	//Even  18 : 1.4020950, 0.4083462
		38 :
			REF <= 32'b0111111001111000_1001001001010110;	//									Odd  19 : 0.9880643, 0.2858130
		39 :
			REF <= 32'b1011001011011011_1100111011110011;	//Even  19 : 1.3973340, 0.4042006
		40 :
			REF <= 32'b0111111000001011_1001000011011100;	//									Odd  20 : 0.9847319, 0.2829308
		41 :
			REF <= 32'b1011001001000001_1100110011011101;	//Even  20 : 1.3926213, 0.4001246
		42 :
			REF <= 32'b0111110110011111_1000111101101000;	//									Odd  21 : 0.9814330, 0.2800968
		43 :
			REF <= 32'b1011000110101000_1100101011001111;	//Even  21 : 1.3879558, 0.3961167
		44 :
			REF <= 32'b0111110100110100_1000110111111011;	//									Odd  22 : 0.9781670, 0.2773098
		45 :
			REF <= 32'b1011000100010001_1100100011001011;	//Even  22 : 1.3833370, 0.3921753
		46 :
			REF <= 32'b0111110011001010_1000110010010100;	//									Odd  23 : 0.9749334, 0.2745687
		47 :
			REF <= 32'b1011000001111011_1100011011001111;	//Even  23 : 1.3787640, 0.3882988
		48 :
			REF <= 32'b0111110001100001_1000101100110010;	//									Odd  24 : 0.9717316, 0.2718725
		49 :
			REF <= 32'b1010111111100110_1100010011011011;	//Even  24 : 1.3742360, 0.3844857
		50 :
			REF <= 32'b0111101111111001_1000100111010111;	//									Odd  25 : 0.9685612, 0.2692201
		51 :
			REF <= 32'b1010111101010100_1100001011101111;	//Even  25 : 1.3697524, 0.3807347
		52 :
			REF <= 32'b0111101110010010_1000100010000001;	//									Odd  26 : 0.9654216, 0.2666105
		53 :
			REF <= 32'b1010111011000010_1100000100001011;	//Even  26 : 1.3653123, 0.3770442
		54 :
			REF <= 32'b0111101100101101_1000011100110000;	//									Odd  27 : 0.9623123, 0.2640428
		55 :
			REF <= 32'b1010111000110010_1011111100101111;	//Even  27 : 1.3609152, 0.3734129
		56 :
			REF <= 32'b0111101011001000_1000010111100101;	//									Odd  28 : 0.9592329, 0.2615161
		57 :
			REF <= 32'b1010110110100011_1011110101011011;	//Even  28 : 1.3565602, 0.3698396
		58 :
			REF <= 32'b0111101001100100_1000010010011111;	//									Odd  29 : 0.9561829, 0.2590294
		59 :
			REF <= 32'b1010110100010110_1011101110001110;	//Even  29 : 1.3522468, 0.3663229
		60 :
			REF <= 32'b0111101000000001_1000001101011110;	//									Odd  30 : 0.9531618, 0.2565819
		61 :
			REF <= 32'b1010110010001010_1011100111001001;	//Even  30 : 1.3479743, 0.3628616
		62 :
			REF <= 32'b0111100110011111_1000001000100010;	//									Odd  31 : 0.9501691, 0.2541727
		63 :
			REF <= 32'b1010101111111111_1011100000001010;	//Even  31 : 1.3437420, 0.3594545
		64 :
			REF <= 32'b0111100100111101_1000000011101100;	//									Odd  32 : 0.9472045, 0.2518010
		65 :
			REF <= 32'b1010101101110110_1011011001010010;	//Even  32 : 1.3395494, 0.3561004
		66 :
			REF <= 32'b0111100011011101_0111111110111001;	//									Odd  33 : 0.9442674, 0.2494659
		67 :
			REF <= 32'b1010101011101110_1011010010100001;	//Even  33 : 1.3353957, 0.3527980
		68 :
			REF <= 32'b0111100001111110_0111111010001100;	//									Odd  34 : 0.9413574, 0.2471667
		69 :
			REF <= 32'b1010101001100111_1011001011110111;	//Even  34 : 1.3312805, 0.3495465
		70 :
			REF <= 32'b0111100000011111_0111110101100011;	//									Odd  35 : 0.9384742, 0.2449026
		71 :
			REF <= 32'b1010100111100001_1011000101010100;	//Even  35 : 1.3272030, 0.3463445
		72 :
			REF <= 32'b0111011111000010_0111110000111111;	//									Odd  36 : 0.9356174, 0.2426728
		73 :
			REF <= 32'b1010100101011101_1010111110110110;	//Even  36 : 1.3231628, 0.3431912
		74 :
			REF <= 32'b0111011101100101_0111101100011111;	//									Odd  37 : 0.9327865, 0.2404767
		75 :
			REF <= 32'b1010100011011010_1010111000011111;	//Even  37 : 1.3191593, 0.3400854
		76 :
			REF <= 32'b0111011100001001_0111101000000100;	//									Odd  38 : 0.9299811, 0.2383135
		77 :
			REF <= 32'b1010100001011000_1010110010001110;	//Even  38 : 1.3151919, 0.3370261
		78 :
			REF <= 32'b0111011010101110_0111100011101100;	//									Odd  39 : 0.9272009, 0.2361825
		79 :
			REF <= 32'b1010011111010111_1010101100000011;	//Even  39 : 1.3112601, 0.3340125
		80 :
			REF <= 32'b0111011001010100_0111011111011001;	//									Odd  40 : 0.9244455, 0.2340831
		81 :
			REF <= 32'b1010011101010111_1010100101111110;	//Even  40 : 1.3073633, 0.3310435
		82 :
			REF <= 32'b0111010111111010_0111011011001010;	//									Odd  41 : 0.9217144, 0.2320147
		83 :
			REF <= 32'b1010011011011001_1010011111111111;	//Even  41 : 1.3035011, 0.3281183
		84 :
			REF <= 32'b0111010110100010_0111010110111111;	//									Odd  42 : 0.9190075, 0.2299765
		85 :
			REF <= 32'b1010011001011011_1010011010000101;	//Even  42 : 1.2996728, 0.3252358
		86 :
			REF <= 32'b0111010101001010_0111010010111000;	//									Odd  43 : 0.9163243, 0.2279679
		87 :
			REF <= 32'b1010010111011111_1010010100010001;	//Even  43 : 1.2958782, 0.3223954
		88 :
			REF <= 32'b0111010011110010_0111001110110100;	//									Odd  44 : 0.9136644, 0.2259885
		89 :
			REF <= 32'b1010010101100100_1010001110100010;	//Even  44 : 1.2921165, 0.3195960
		90 :
			REF <= 32'b0111010010011100_0111001010110101;	//									Odd  45 : 0.9110276, 0.2240375
		91 :
			REF <= 32'b1010010011101001_1010001000111000;	//Even  45 : 1.2883875, 0.3168369
		92 :
			REF <= 32'b0111010001000110_0111000110111000;	//									Odd  46 : 0.9084134, 0.2221144
		93 :
			REF <= 32'b1010010001110000_1010000011010011;	//Even  46 : 1.2846905, 0.3141173
		94 :
			REF <= 32'b0111001111110001_0111000011000000;	//									Odd  47 : 0.9058216, 0.2202187
		95 :
			REF <= 32'b1010001111111000_1001111101110100;	//Even  47 : 1.2810252, 0.3114363
		96 :
			REF <= 32'b0111001110011101_0110111111001011;	//									Odd  48 : 0.9032519, 0.2183498
		97 :
			REF <= 32'b1010001110000001_1001111000011010;	//Even  48 : 1.2773911, 0.3087933
		98 :
			REF <= 32'b0111001101001010_0110111011011010;	//									Odd  49 : 0.9007040, 0.2165072
		99 :
			REF <= 32'b1010001100001011_1001110011000100;	//Even  49 : 1.2737877, 0.3061875
		100 :
			REF <= 32'b0111001011110111_0110110111101011;	//									Odd  50 : 0.8981774, 0.2146904
		101 :
			REF <= 32'b1010001010010110_1001101101110011;	//Even  50 : 1.2702147, 0.3036181
		102 :
			REF <= 32'b0111001010100101_0110110100000001;	//									Odd  51 : 0.8956720, 0.2128988
		103 :
			REF <= 32'b1010001000100010_1001101000100111;	//Even  51 : 1.2666715, 0.3010844
		104 :
			REF <= 32'b0111001001010011_0110110000011001;	//									Odd  52 : 0.8931875, 0.2111320
		105 :
			REF <= 32'b1010000110101111_1001100011100000;	//Even  52 : 1.2631578, 0.2985858
		106 :
			REF <= 32'b0111001000000011_0110101100110101;	//									Odd  53 : 0.8907235, 0.2093896
		107 :
			REF <= 32'b1010000100111100_1001011110011101;	//Even  53 : 1.2596734, 0.2961215
		108 :
			REF <= 32'b0111000110110011_0110101001010011;	//									Odd  54 : 0.8882799, 0.2076709
		109 :
			REF <= 32'b1010000011001011_1001011001011110;	//Even  54 : 1.2562174, 0.2936910
		110 :
			REF <= 32'b0111000101100011_0110100101110101;	//									Odd  55 : 0.8858562, 0.2059756
		111 :
			REF <= 32'b1010000001011011_1001010100100100;	//Even  55 : 1.2527899, 0.2912935
		112 :
			REF <= 32'b0111000100010100_0110100010011010;	//									Odd  56 : 0.8834522, 0.2043033
		113 :
			REF <= 32'b1001111111101100_1001001111101110;	//Even  56 : 1.2493901, 0.2889285
		114 :
			REF <= 32'b0111000011000110_0110011111000010;	//									Odd  57 : 0.8810677, 0.2026535
		115 :
			REF <= 32'b1001111101111101_1001001010111100;	//Even  57 : 1.2460179, 0.2865953
		116 :
			REF <= 32'b0111000001111001_0110011011101100;	//									Odd  58 : 0.8787024, 0.2010258
		117 :
			REF <= 32'b1001111100001111_1001000110001110;	//Even  58 : 1.2426729, 0.2842934
		118 :
			REF <= 32'b0111000000101100_0110011000011010;	//									Odd  59 : 0.8763561, 0.1994197
		119 :
			REF <= 32'b1001111010100011_1001000001100101;	//Even  59 : 1.2393547, 0.2820220
		120 :
			REF <= 32'b0110111111100000_0110010101001010;	//									Odd  60 : 0.8740284, 0.1978349
		121 :
			REF <= 32'b1001111000110111_1000111100111111;	//Even  60 : 1.2360629, 0.2797808
		122 :
			REF <= 32'b0110111110010100_0110010001111101;	//									Odd  61 : 0.8717192, 0.1962710
		123 :
			REF <= 32'b1001110111001100_1000111000011101;	//Even  61 : 1.2327971, 0.2775691
		124 :
			REF <= 32'b0110111101001001_0110001110110011;	//									Odd  62 : 0.8694283, 0.1947276
		125 :
			REF <= 32'b1001110101100010_1000110011111111;	//Even  62 : 1.2295573, 0.2753864
		126 :
			REF <= 32'b0110111011111110_0110001011101011;	//									Odd  63 : 0.8671553, 0.1932043
		127 :
			REF <= 32'b1001110011111000_1000101111100101;	//Even  63 : 1.2263427, 0.2732321
		128 :
			REF <= 32'b0110111010110101_0110001000100110;	//									Odd  64 : 0.8649000, 0.1917008
		129 :
			REF <= 32'b1001110010010000_1000101011001110;	//Even  64 : 1.2231532, 0.2711058
		130 :
			REF <= 32'b0110111001101011_0110000101100100;	//									Odd  65 : 0.8626622, 0.1902166
		131 :
			REF <= 32'b1001110000101000_1000100110111011;	//Even  65 : 1.2199886, 0.2690070
		132 :
			REF <= 32'b0110111000100010_0110000010100100;	//									Odd  66 : 0.8604417, 0.1887516
		133 :
			REF <= 32'b1001101111000001_1000100010101011;	//Even  66 : 1.2168483, 0.2669350
		134 :
			REF <= 32'b0110110111011010_0101111111100110;	//									Odd  67 : 0.8582382, 0.1873052
		135 :
			REF <= 32'b1001101101011011_1000011110011111;	//Even  67 : 1.2137321, 0.2648895
		136 :
			REF <= 32'b0110110110010011_0101111100101011;	//									Odd  68 : 0.8560516, 0.1858772
		137 :
			REF <= 32'b1001101011110110_1000011010010110;	//Even  68 : 1.2106398, 0.2628701
		138 :
			REF <= 32'b0110110101001011_0101111001110010;	//									Odd  69 : 0.8538817, 0.1844673
		139 :
			REF <= 32'b1001101010010001_1000010110010001;	//Even  69 : 1.2075710, 0.2608761
		140 :
			REF <= 32'b0110110100000101_0101110110111100;	//									Odd  70 : 0.8517281, 0.1830751
		141 :
			REF <= 32'b1001101000101101_1000010010001111;	//Even  70 : 1.2045255, 0.2589072
		142 :
			REF <= 32'b0110110010111111_0101110100000111;	//									Odd  71 : 0.8495908, 0.1817003
		143 :
			REF <= 32'b1001100111001010_1000001110010000;	//Even  71 : 1.2015028, 0.2569630
		144 :
			REF <= 32'b0110110001111001_0101110001010101;	//									Odd  72 : 0.8474694, 0.1803426
		145 :
			REF <= 32'b1001100101101000_1000001010010100;	//Even  72 : 1.1985028, 0.2550430
		146 :
			REF <= 32'b0110110000110100_0101101110100110;	//									Odd  73 : 0.8453639, 0.1790018
		147 :
			REF <= 32'b1001100100000110_1000000110011100;	//Even  73 : 1.1955252, 0.2531468
		148 :
			REF <= 32'b0110101111110000_0101101011111000;	//									Odd  74 : 0.8432741, 0.1776775
		149 :
			REF <= 32'b1001100010100110_1000000010100110;	//Even  74 : 1.1925696, 0.2512739
		150 :
			REF <= 32'b0110101110101100_0101101001001101;	//									Odd  75 : 0.8411996, 0.1763694
		151 :
			REF <= 32'b1001100001000101_0111111110110100;	//Even  75 : 1.1896359, 0.2494241
		152 :
			REF <= 32'b0110101101101000_0101100110100011;	//									Odd  76 : 0.8391403, 0.1750774
		153 :
			REF <= 32'b1001011111100110_0111111011000101;	//Even  76 : 1.1867236, 0.2475968
		154 :
			REF <= 32'b0110101100100101_0101100011111100;	//									Odd  77 : 0.8370962, 0.1738010
		155 :
			REF <= 32'b1001011110000111_0111110111011000;	//Even  77 : 1.1838326, 0.2457917
		156 :
			REF <= 32'b0110101011100011_0101100001010111;	//									Odd  78 : 0.8350668, 0.1725400
		157 :
			REF <= 32'b1001011100101001_0111110011101110;	//Even  78 : 1.1809628, 0.2440085
		158 :
			REF <= 32'b0110101010100001_0101011110110011;	//									Odd  79 : 0.8330522, 0.1712943
		159 :
			REF <= 32'b1001011011001100_0111110000000111;	//Even  79 : 1.1781137, 0.2422467
		160 :
			REF <= 32'b0110101001011111_0101011100010010;	//									Odd  80 : 0.8310520, 0.1700634
		161 :
			REF <= 32'b1001011001101111_0111101100100011;	//Even  80 : 1.1752851, 0.2405060
		162 :
			REF <= 32'b0110101000011110_0101011001110011;	//									Odd  81 : 0.8290662, 0.1688472
		163 :
			REF <= 32'b1001011000010011_0111101001000010;	//Even  81 : 1.1724768, 0.2387860
		164 :
			REF <= 32'b0110100111011110_0101010111010101;	//									Odd  82 : 0.8270946, 0.1676455
		165 :
			REF <= 32'b1001010110111000_0111100101100011;	//Even  82 : 1.1696885, 0.2370865
		166 :
			REF <= 32'b0110100110011110_0101010100111001;	//									Odd  83 : 0.8251370, 0.1664579
		167 :
			REF <= 32'b1001010101011101_0111100010000111;	//Even  83 : 1.1669199, 0.2354070
		168 :
			REF <= 32'b0110100101011110_0101010010100000;	//									Odd  84 : 0.8231932, 0.1652843
		169 :
			REF <= 32'b1001010100000011_0111011110101101;	//Even  84 : 1.1641710, 0.2337473
		170 :
			REF <= 32'b0110100100011111_0101010000001000;	//									Odd  85 : 0.8212631, 0.1641244
		171 :
			REF <= 32'b1001010010101010_0111011011010110;	//Even  85 : 1.1614414, 0.2321070
		172 :
			REF <= 32'b0110100011100000_0101001101110001;	//									Odd  86 : 0.8193465, 0.1629780
		173 :
			REF <= 32'b1001010001010001_0111011000000010;	//Even  86 : 1.1587309, 0.2304857
		174 :
			REF <= 32'b0110100010100001_0101001011011101;	//									Odd  87 : 0.8174433, 0.1618449
		175 :
			REF <= 32'b1001001111111001_0111010100110000;	//Even  87 : 1.1560394, 0.2288833
		176 :
			REF <= 32'b0110100001100100_0101001001001010;	//									Odd  88 : 0.8155532, 0.1607249
		177 :
			REF <= 32'b1001001110100001_0111010001100000;	//Even  88 : 1.1533664, 0.2272993
		178 :
			REF <= 32'b0110100000100110_0101000110111001;	//									Odd  89 : 0.8136762, 0.1596177
		179 :
			REF <= 32'b1001001101001010_0111001110010011;	//Even  89 : 1.1507119, 0.2257335
		180 :
			REF <= 32'b0110011111101001_0101000100101001;	//									Odd  90 : 0.8118121, 0.1585232
		181 :
			REF <= 32'b1001001011110100_0111001011001000;	//Even  90 : 1.1480757, 0.2241856
		182 :
			REF <= 32'b0110011110101100_0101000010011100;	//									Odd  91 : 0.8099608, 0.1574411
		183 :
			REF <= 32'b1001001010011110_0111000111111111;	//Even  91 : 1.1454575, 0.2226554
		184 :
			REF <= 32'b0110011101110000_0101000000001111;	//									Odd  92 : 0.8081220, 0.1563713
		185 :
			REF <= 32'b1001001001001001_0111000100111001;	//Even  92 : 1.1428572, 0.2211424
		186 :
			REF <= 32'b0110011100110100_0100111110000101;	//									Odd  93 : 0.8062958, 0.1553136
		187 :
			REF <= 32'b1001000111110100_0111000001110101;	//Even  93 : 1.1402744, 0.2196465
		188 :
			REF <= 32'b0110011011111001_0100111011111100;	//									Odd  94 : 0.8044818, 0.1542677
		189 :
			REF <= 32'b1001000110100000_0110111110110011;	//Even  94 : 1.1377091, 0.2181674
		190 :
			REF <= 32'b0110011010111110_0100111001110100;	//									Odd  95 : 0.8026801, 0.1532335
		191 :
			REF <= 32'b1001000101001100_0110111011110011;	//Even  95 : 1.1351610, 0.2167049
		192 :
			REF <= 32'b0110011010000011_0100110111101110;	//									Odd  96 : 0.8008904, 0.1522108
		193 :
			REF <= 32'b1001000011111010_0110111000110110;	//Even  96 : 1.1326300, 0.2152586
		194 :
			REF <= 32'b0110011001001001_0100110101101010;	//									Odd  97 : 0.7991126, 0.1511994
		195 :
			REF <= 32'b1001000010100111_0110110101111010;	//Even  97 : 1.1301159, 0.2138283
		196 :
			REF <= 32'b0110011000001111_0100110011100110;	//									Odd  98 : 0.7973466, 0.1501992
		197 :
			REF <= 32'b1001000001010101_0110110011000001;	//Even  98 : 1.1276183, 0.2124138
		198 :
			REF <= 32'b0110010111010101_0100110001100101;	//									Odd  99 : 0.7955922, 0.1492100
		199 :
			REF <= 32'b1001000000000100_0110110000001010;	//Even  99 : 1.1251373, 0.2110148
		200 :
			REF <= 32'b0110010110011100_0100101111100101;	//									Odd 100 : 0.7938495, 0.1482316
		201 :
			REF <= 32'b1000111110110011_0110101101010100;	//Even 100 : 1.1226727, 0.2096311
		202 :
			REF <= 32'b0110010101100100_0100101101100110;	//									Odd 101 : 0.7921180, 0.1472638
		203 :
			REF <= 32'b1000111101100011_0110101010100001;	//Even 101 : 1.1202241, 0.2082624
		204 :
			REF <= 32'b0110010100101011_0100101011101000;	//									Odd 102 : 0.7903979, 0.1463065
		205 :
			REF <= 32'b1000111100010011_0110100111101111;	//Even 102 : 1.1177914, 0.2069086
		206 :
			REF <= 32'b0110010011110011_0100101001101100;	//									Odd 103 : 0.7886890, 0.1453595
		207 :
			REF <= 32'b1000111011000100_0110100101000000;	//Even 103 : 1.1153746, 0.2055694
		208 :
			REF <= 32'b0110010010111100_0100100111110001;	//									Odd 104 : 0.7869910, 0.1444227
		209 :
			REF <= 32'b1000111001110101_0110100010010010;	//Even 104 : 1.1129733, 0.2042446
		210 :
			REF <= 32'b0110010010000100_0100100101111000;	//									Odd 105 : 0.7853040, 0.1434959
		211 :
			REF <= 32'b1000111000100111_0110011111100110;	//Even 105 : 1.1105876, 0.2029339
		212 :
			REF <= 32'b0110010001001101_0100100100000000;	//									Odd 106 : 0.7836277, 0.1425790
		213 :
			REF <= 32'b1000110111011010_0110011100111100;	//Even 106 : 1.1082170, 0.2016372
		214 :
			REF <= 32'b0110010000010111_0100100010001001;	//									Odd 107 : 0.7819623, 0.1416719
		215 :
			REF <= 32'b1000110110001100_0110011010010100;	//Even 107 : 1.1058617, 0.2003543
		216 :
			REF <= 32'b0110001111100001_0100100000010011;	//									Odd 108 : 0.7803073, 0.1407743
		217 :
			REF <= 32'b1000110101000000_0110010111101110;	//Even 108 : 1.1035212, 0.1990849
		218 :
			REF <= 32'b0110001110101011_0100011110011111;	//									Odd 109 : 0.7786628, 0.1398861
		219 :
			REF <= 32'b1000110011110011_0110010101001001;	//Even 109 : 1.1011956, 0.1978288
		220 :
			REF <= 32'b0110001101110101_0100011100101011;	//									Odd 110 : 0.7770287, 0.1390072
		221 :
			REF <= 32'b1000110010101000_0110010010100110;	//Even 110 : 1.0988845, 0.1965859
		222 :
			REF <= 32'b0110001101000000_0100011010111001;	//									Odd 111 : 0.7754048, 0.1381375
		223 :
			REF <= 32'b1000110001011100_0110010000000101;	//Even 111 : 1.0965880, 0.1953560
		224 :
			REF <= 32'b0110001100001011_0100011001001001;	//									Odd 112 : 0.7737911, 0.1372769
		225 :
			REF <= 32'b1000110000010010_0110001101100110;	//Even 112 : 1.0943058, 0.1941388
		226 :
			REF <= 32'b0110001011010111_0100010111011001;	//									Odd 113 : 0.7721874, 0.1364251
		227 :
			REF <= 32'b1000101111000111_0110001011001000;	//Even 113 : 1.0920378, 0.1929342
		228 :
			REF <= 32'b0110001010100010_0100010101101011;	//									Odd 114 : 0.7705936, 0.1355821
		229 :
			REF <= 32'b1000101101111110_0110001000101100;	//Even 114 : 1.0897839, 0.1917420
		230 :
			REF <= 32'b0110001001101110_0100010011111101;	//									Odd 115 : 0.7690096, 0.1347477
		231 :
			REF <= 32'b1000101100110100_0110000110010001;	//Even 115 : 1.0875438, 0.1905621
		232 :
			REF <= 32'b0110001000111011_0100010010010001;	//									Odd 116 : 0.7674354, 0.1339219
		233 :
			REF <= 32'b1000101011101011_0110000011111000;	//Even 116 : 1.0853175, 0.1893942
		234 :
			REF <= 32'b0110001000001000_0100010000100110;	//									Odd 117 : 0.7658707, 0.1331045
		235 :
			REF <= 32'b1000101010100011_0110000001100000;	//Even 117 : 1.0831048, 0.1882382
		236 :
			REF <= 32'b0110000111010101_0100001110111100;	//									Odd 118 : 0.7643157, 0.1322954
		237 :
			REF <= 32'b1000101001011011_0101111111001010;	//Even 118 : 1.0809057, 0.1870939
		238 :
			REF <= 32'b0110000110100010_0100001101010011;	//									Odd 119 : 0.7627701, 0.1314944
		239 :
			REF <= 32'b1000101000010011_0101111100110110;	//Even 119 : 1.0787197, 0.1859611
		240 :
			REF <= 32'b0110000101110000_0100001011101011;	//									Odd 120 : 0.7612337, 0.1307014
		241 :
			REF <= 32'b1000100111001100_0101111010100011;	//Even 120 : 1.0765471, 0.1848398
		242 :
			REF <= 32'b0110000100111110_0100001010000100;	//									Odd 121 : 0.7597067, 0.1299164
		243 :
			REF <= 32'b1000100110000101_0101111000010001;	//Even 121 : 1.0743876, 0.1837296
		244 :
			REF <= 32'b0110000100001100_0100001000011110;	//									Odd 122 : 0.7581888, 0.1291393
		245 :
			REF <= 32'b1000100100111111_0101110110000001;	//Even 122 : 1.0722409, 0.1826305
		246 :
			REF <= 32'b0110000011011010_0100000110111001;	//									Odd 123 : 0.7566800, 0.1283698
		247 :
			REF <= 32'b1000100011111001_0101110011110011;	//Even 123 : 1.0701071, 0.1815424
		248 :
			REF <= 32'b0110000010101001_0100000101010101;	//									Odd 124 : 0.7551801, 0.1276080
		249 :
			REF <= 32'b1000100010110011_0101110001100101;	//Even 124 : 1.0679860, 0.1804650
		250 :
			REF <= 32'b0110000001111000_0100000011110010;	//									Odd 125 : 0.7536892, 0.1268537
		251 :
			REF <= 32'b1000100001101110_0101101111011010;	//Even 125 : 1.0658774, 0.1793982
		252 :
			REF <= 32'b0110000001001000_0100000010010001;	//									Odd 126 : 0.7522070, 0.1261067
		253 :
			REF <= 32'b1000100000101001_0101101101001111;	//Even 126 : 1.0637813, 0.1783419
		254 :
			REF <= 32'b0110000000011000_0100000000110000;	//									Odd 127 : 0.7507335, 0.1253671
		255 :
			REF <= 32'b1000011111100101_0101101011000110;	//Even 127 : 1.0616975, 0.1772959
	endcase
end

endmodule
