//================================================================================
// Copyright (c) 2013 ~ 2019. HyungKi Jeong(clonextop@gmail.com)
// All rights reserved.
// 
// The 3-Clause BSD License (https://opensource.org/licenses/BSD-3-Clause)
// 
// Redistribution and use in source and binary forms,
// with or without modification, are permitted provided
// that the following conditions are met:
// 
// 1. Redistributions of source code must retain the above copyright notice,
//    this list of conditions and the following disclaimer.
// 
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
// 
// 3. Neither the name of the copyright holder nor the names of its contributors
//    may be used to endorse or promote products derived from this software
//    without specific prior written permission.
// 
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
// THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
// PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS
// BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE
// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
// HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
// STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN
// ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY
// OF SUCH DAMAGE.
// 
// Title : Meitner processor v1.1
// Rev.  : 10/31/2019 Thu (clonextop@gmail.com)
//================================================================================
`include "MTSP_Defines.vh"

module MTSP_SF_RCP_LUT(CLK, index, REF);
// port definition -----------------------------------------------------------
input	CLK;
input	[7:0]		index;		// LUT index
output reg	[22:0]	REF;		// Reference Value

// register definition & assignment ------------------------------------------

// behavior code -------------------------------------------------------------
`ALWAYS_CLOCK begin
	case(index) //	  Reference     Reference^2
		0 :
			REF <= 23'b1111111_1111111100000000;	// 2
		1 :
			REF <= 23'b1111101_1111110100000010;	// 2
		2 :
			REF <= 23'b1111011_1111101100000110;	// 2
		3 :
			REF <= 23'b1111001_1111100100001100;	// 2
		4 :
			REF <= 23'b1110111_1111011100010100;	// 2
		5 :
			REF <= 23'b1110101_1111010100011110;	// 2
		6 :
			REF <= 23'b1110011_1111001100101010;	// 2
		7 :
			REF <= 23'b1110001_1111000100111000;	// 1
		8 :
			REF <= 23'b1110000_1111000001000000;	// 2
		9 :
			REF <= 23'b1101110_1110111001010001;	// 2
		10 :
			REF <= 23'b1101100_1110110001100100;	// 2
		11 :
			REF <= 23'b1101010_1110101001111001;	// 2
		12 :
			REF <= 23'b1101000_1110100010010000;	// 2
		13 :
			REF <= 23'b1100110_1110011010101001;	// 1
		14 :
			REF <= 23'b1100101_1110010110110110;	// 2
		15 :
			REF <= 23'b1100011_1110001111010010;	// 2
		16 :
			REF <= 23'b1100001_1110000111110000;	// 2
		17 :
			REF <= 23'b1011111_1110000000010000;	// 2
		18 :
			REF <= 23'b1011101_1101111000110010;	// 1
		19 :
			REF <= 23'b1011100_1101110101000100;	// 2
		20 :
			REF <= 23'b1011010_1101101101101001;	// 2
		21 :
			REF <= 23'b1011000_1101100110010000;	// 1
		22 :
			REF <= 23'b1010111_1101100010100100;	// 2
		23 :
			REF <= 23'b1010101_1101011011001110;	// 2
		24 :
			REF <= 23'b1010011_1101010011111010;	// 1
		25 :
			REF <= 23'b1010010_1101010000010001;	// 2
		26 :
			REF <= 23'b1010000_1101001001000000;	// 2
		27 :
			REF <= 23'b1001110_1101000001110001;	// 1
		28 :
			REF <= 23'b1001101_1100111110001010;	// 2
		29 :
			REF <= 23'b1001011_1100110110111110;	// 2
		30 :
			REF <= 23'b1001001_1100101111110100;	// 1
		31 :
			REF <= 23'b1001000_1100101100010000;	// 2
		32 :
			REF <= 23'b1000110_1100100101001001;	// 1
		33 :
			REF <= 23'b1000101_1100100001100110;	// 2
		34 :
			REF <= 23'b1000011_1100011010100010;	// 1
		35 :
			REF <= 23'b1000010_1100010111000001;	// 2
		36 :
			REF <= 23'b1000000_1100010000000000;	// 1
		37 :
			REF <= 23'b0111111_1100001100100000;	// 2
		38 :
			REF <= 23'b0111101_1100000101100010;	// 1
		39 :
			REF <= 23'b0111100_1100000010000100;	// 2
		40 :
			REF <= 23'b0111010_1011111011001001;	// 1
		41 :
			REF <= 23'b0111001_1011110111101100;	// 2
		42 :
			REF <= 23'b0110111_1011110000110100;	// 1
		43 :
			REF <= 23'b0110110_1011101101011001;	// 2
		44 :
			REF <= 23'b0110100_1011100110100100;	// 1
		45 :
			REF <= 23'b0110011_1011100011001010;	// 2
		46 :
			REF <= 23'b0110001_1011011100011000;	// 1
		47 :
			REF <= 23'b0110000_1011011001000000;	// 2
		48 :
			REF <= 23'b0101110_1011010010010001;	// 1
		49 :
			REF <= 23'b0101101_1011001110111010;	// 1
		50 :
			REF <= 23'b0101100_1011001011100100;	// 2
		51 :
			REF <= 23'b0101010_1011000100111001;	// 1
		52 :
			REF <= 23'b0101001_1011000001100100;	// 2
		53 :
			REF <= 23'b0100111_1010111010111100;	// 1
		54 :
			REF <= 23'b0100110_1010110111101001;	// 1
		55 :
			REF <= 23'b0100101_1010110100010110;	// 2
		56 :
			REF <= 23'b0100011_1010101101110010;	// 1
		57 :
			REF <= 23'b0100010_1010101010100001;	// 1
		58 :
			REF <= 23'b0100001_1010100111010000;	// 2
		59 :
			REF <= 23'b0011111_1010100000110000;	// 1
		60 :
			REF <= 23'b0011110_1010011101100001;	// 1
		61 :
			REF <= 23'b0011101_1010011010010010;	// 1
		62 :
			REF <= 23'b0011100_1010010111000100;	// 2
		63 :
			REF <= 23'b0011010_1010010000101001;	// 1
		64 :
			REF <= 23'b0011001_1010001101011100;	// 1
		65 :
			REF <= 23'b0011000_1010001010010000;	// 2
		66 :
			REF <= 23'b0010110_1010000011111001;	// 1
		67 :
			REF <= 23'b0010101_1010000000101110;	// 1
		68 :
			REF <= 23'b0010100_1001111101100100;	// 1
		69 :
			REF <= 23'b0010011_1001111010011010;	// 2
		70 :
			REF <= 23'b0010001_1001110100001000;	// 1
		71 :
			REF <= 23'b0010000_1001110001000000;	// 1
		72 :
			REF <= 23'b0001111_1001101101111000;	// 1
		73 :
			REF <= 23'b0001110_1001101010110001;	// 1
		74 :
			REF <= 23'b0001101_1001100111101010;	// 2
		75 :
			REF <= 23'b0001011_1001100001011110;	// 1
		76 :
			REF <= 23'b0001010_1001011110011001;	// 1
		77 :
			REF <= 23'b0001001_1001011011010100;	// 1
		78 :
			REF <= 23'b0001000_1001011000010000;	// 1
		79 :
			REF <= 23'b0000111_1001010101001100;	// 1
		80 :
			REF <= 23'b0000110_1001010010001001;	// 2
		81 :
			REF <= 23'b0000100_1001001100000100;	// 1
		82 :
			REF <= 23'b0000011_1001001001000010;	// 1
		83 :
			REF <= 23'b0000010_1001000110000001;	// 1
		84 :
			REF <= 23'b0000001_1001000011000000;	// 1
		85 :
			REF <= 23'b0000000_1001000000000000;	// 1
		86 :
			REF <= 23'b1111111_1000111101000000;	// 1
		87 :
			REF <= 23'b1111110_1000111010000001;	// 2
		88 :
			REF <= 23'b1111100_1000110100000100;	// 1
		89 :
			REF <= 23'b1111011_1000110001000110;	// 1
		90 :
			REF <= 23'b1111010_1000101110001001;	// 1
		91 :
			REF <= 23'b1111001_1000101011001100;	// 1
		92 :
			REF <= 23'b1111000_1000101000010000;	// 1
		93 :
			REF <= 23'b1110111_1000100101010100;	// 1
		94 :
			REF <= 23'b1110110_1000100010011001;	// 1
		95 :
			REF <= 23'b1110101_1000011111011110;	// 1
		96 :
			REF <= 23'b1110100_1000011100100100;	// 1
		97 :
			REF <= 23'b1110011_1000011001101010;	// 1
		98 :
			REF <= 23'b1110010_1000010110110001;	// 1
		99 :
			REF <= 23'b1110001_1000010011111000;	// 1
		100 :
			REF <= 23'b1110000_1000010001000000;	// 1
		101 :
			REF <= 23'b1101111_1000001110001000;	// 1
		102 :
			REF <= 23'b1101110_1000001011010001;	// 1
		103 :
			REF <= 23'b1101101_1000001000011010;	// 1
		104 :
			REF <= 23'b1101100_1000000101100100;	// 1
		105 :
			REF <= 23'b1101011_1000000010101110;	// 1
		106 :
			REF <= 23'b1101010_0111111111111001;	// 1
		107 :
			REF <= 23'b1101001_0111111101000100;	// 1
		108 :
			REF <= 23'b1101000_0111111010010000;	// 1
		109 :
			REF <= 23'b1100111_0111110111011100;	// 1
		110 :
			REF <= 23'b1100110_0111110100101001;	// 1
		111 :
			REF <= 23'b1100101_0111110001110110;	// 1
		112 :
			REF <= 23'b1100100_0111101111000100;	// 1
		113 :
			REF <= 23'b1100011_0111101100010010;	// 1
		114 :
			REF <= 23'b1100010_0111101001100001;	// 1
		115 :
			REF <= 23'b1100001_0111100110110000;	// 1
		116 :
			REF <= 23'b1100000_0111100100000000;	// 1
		117 :
			REF <= 23'b1011111_0111100001010000;	// 1
		118 :
			REF <= 23'b1011110_0111011110100001;	// 1
		119 :
			REF <= 23'b1011101_0111011011110010;	// 1
		120 :
			REF <= 23'b1011100_0111011001000100;	// 1
		121 :
			REF <= 23'b1011011_0111010110010110;	// 1
		122 :
			REF <= 23'b1011010_0111010011101001;	// 1
		123 :
			REF <= 23'b1011001_0111010000111100;	// 1
		124 :
			REF <= 23'b1011000_0111001110010000;	// 0
		125 :
			REF <= 23'b1011000_0111001110010000;	// 1
		126 :
			REF <= 23'b1010111_0111001011100100;	// 1
		127 :
			REF <= 23'b1010110_0111001000111001;	// 1
		128 :
			REF <= 23'b1010101_0111000110001110;	// 1
		129 :
			REF <= 23'b1010100_0111000011100100;	// 1
		130 :
			REF <= 23'b1010011_0111000000111010;	// 1
		131 :
			REF <= 23'b1010010_0110111110010001;	// 1
		132 :
			REF <= 23'b1010001_0110111011101000;	// 0
		133 :
			REF <= 23'b1010001_0110111011101000;	// 1
		134 :
			REF <= 23'b1010000_0110111001000000;	// 1
		135 :
			REF <= 23'b1001111_0110110110011000;	// 1
		136 :
			REF <= 23'b1001110_0110110011110001;	// 1
		137 :
			REF <= 23'b1001101_0110110001001010;	// 1
		138 :
			REF <= 23'b1001100_0110101110100100;	// 1
		139 :
			REF <= 23'b1001011_0110101011111110;	// 0
		140 :
			REF <= 23'b1001011_0110101011111110;	// 1
		141 :
			REF <= 23'b1001010_0110101001011001;	// 1
		142 :
			REF <= 23'b1001001_0110100110110100;	// 1
		143 :
			REF <= 23'b1001000_0110100100010000;	// 1
		144 :
			REF <= 23'b1000111_0110100001101100;	// 1
		145 :
			REF <= 23'b1000110_0110011111001001;	// 0
		146 :
			REF <= 23'b1000110_0110011111001001;	// 1
		147 :
			REF <= 23'b1000101_0110011100100110;	// 1
		148 :
			REF <= 23'b1000100_0110011010000100;	// 1
		149 :
			REF <= 23'b1000011_0110010111100010;	// 1
		150 :
			REF <= 23'b1000010_0110010101000001;	// 0
		151 :
			REF <= 23'b1000010_0110010101000001;	// 1
		152 :
			REF <= 23'b1000001_0110010010100000;	// 1
		153 :
			REF <= 23'b1000000_0110010000000000;	// 1
		154 :
			REF <= 23'b0111111_0110001101100000;	// 0
		155 :
			REF <= 23'b0111111_0110001101100000;	// 1
		156 :
			REF <= 23'b0111110_0110001011000001;	// 1
		157 :
			REF <= 23'b0111101_0110001000100010;	// 1
		158 :
			REF <= 23'b0111100_0110000110000100;	// 1
		159 :
			REF <= 23'b0111011_0110000011100110;	// 0
		160 :
			REF <= 23'b0111011_0110000011100110;	// 1
		161 :
			REF <= 23'b0111010_0110000001001001;	// 1
		162 :
			REF <= 23'b0111001_0101111110101100;	// 1
		163 :
			REF <= 23'b0111000_0101111100010000;	// 0
		164 :
			REF <= 23'b0111000_0101111100010000;	// 1
		165 :
			REF <= 23'b0110111_0101111001110100;	// 1
		166 :
			REF <= 23'b0110110_0101110111011001;	// 1
		167 :
			REF <= 23'b0110101_0101110100111110;	// 0
		168 :
			REF <= 23'b0110101_0101110100111110;	// 1
		169 :
			REF <= 23'b0110100_0101110010100100;	// 1
		170 :
			REF <= 23'b0110011_0101110000001010;	// 0
		171 :
			REF <= 23'b0110011_0101110000001010;	// 1
		172 :
			REF <= 23'b0110010_0101101101110001;	// 1
		173 :
			REF <= 23'b0110001_0101101011011000;	// 1
		174 :
			REF <= 23'b0110000_0101101001000000;	// 0
		175 :
			REF <= 23'b0110000_0101101001000000;	// 1
		176 :
			REF <= 23'b0101111_0101100110101000;	// 1
		177 :
			REF <= 23'b0101110_0101100100010001;	// 0
		178 :
			REF <= 23'b0101110_0101100100010001;	// 1
		179 :
			REF <= 23'b0101101_0101100001111010;	// 1
		180 :
			REF <= 23'b0101100_0101011111100100;	// 0
		181 :
			REF <= 23'b0101100_0101011111100100;	// 1
		182 :
			REF <= 23'b0101011_0101011101001110;	// 1
		183 :
			REF <= 23'b0101010_0101011010111001;	// 0
		184 :
			REF <= 23'b0101010_0101011010111001;	// 1
		185 :
			REF <= 23'b0101001_0101011000100100;	// 1
		186 :
			REF <= 23'b0101000_0101010110010000;	// 0
		187 :
			REF <= 23'b0101000_0101010110010000;	// 1
		188 :
			REF <= 23'b0100111_0101010011111100;	// 1
		189 :
			REF <= 23'b0100110_0101010001101001;	// 0
		190 :
			REF <= 23'b0100110_0101010001101001;	// 1
		191 :
			REF <= 23'b0100101_0101001111010110;	// 1
		192 :
			REF <= 23'b0100100_0101001101000100;	// 0
		193 :
			REF <= 23'b0100100_0101001101000100;	// 1
		194 :
			REF <= 23'b0100011_0101001010110010;	// 1
		195 :
			REF <= 23'b0100010_0101001000100001;	// 0
		196 :
			REF <= 23'b0100010_0101001000100001;	// 1
		197 :
			REF <= 23'b0100001_0101000110010000;	// 1
		198 :
			REF <= 23'b0100000_0101000100000000;	// 0
		199 :
			REF <= 23'b0100000_0101000100000000;	// 1
		200 :
			REF <= 23'b0011111_0101000001110000;	// 1
		201 :
			REF <= 23'b0011110_0100111111100001;	// 0
		202 :
			REF <= 23'b0011110_0100111111100001;	// 1
		203 :
			REF <= 23'b0011101_0100111101010010;	// 0
		204 :
			REF <= 23'b0011101_0100111101010010;	// 1
		205 :
			REF <= 23'b0011100_0100111011000100;	// 1
		206 :
			REF <= 23'b0011011_0100111000110110;	// 0
		207 :
			REF <= 23'b0011011_0100111000110110;	// 1
		208 :
			REF <= 23'b0011010_0100110110101001;	// 0
		209 :
			REF <= 23'b0011010_0100110110101001;	// 1
		210 :
			REF <= 23'b0011001_0100110100011100;	// 1
		211 :
			REF <= 23'b0011000_0100110010010000;	// 0
		212 :
			REF <= 23'b0011000_0100110010010000;	// 1
		213 :
			REF <= 23'b0010111_0100110000000100;	// 0
		214 :
			REF <= 23'b0010111_0100110000000100;	// 1
		215 :
			REF <= 23'b0010110_0100101101111001;	// 1
		216 :
			REF <= 23'b0010101_0100101011101110;	// 0
		217 :
			REF <= 23'b0010101_0100101011101110;	// 1
		218 :
			REF <= 23'b0010100_0100101001100100;	// 0
		219 :
			REF <= 23'b0010100_0100101001100100;	// 1
		220 :
			REF <= 23'b0010011_0100100111011010;	// 1
		221 :
			REF <= 23'b0010010_0100100101010001;	// 0
		222 :
			REF <= 23'b0010010_0100100101010001;	// 1
		223 :
			REF <= 23'b0010001_0100100011001000;	// 0
		224 :
			REF <= 23'b0010001_0100100011001000;	// 1
		225 :
			REF <= 23'b0010000_0100100001000000;	// 0
		226 :
			REF <= 23'b0010000_0100100001000000;	// 1
		227 :
			REF <= 23'b0001111_0100011110111000;	// 0
		228 :
			REF <= 23'b0001111_0100011110111000;	// 1
		229 :
			REF <= 23'b0001110_0100011100110001;	// 1
		230 :
			REF <= 23'b0001101_0100011010101010;	// 0
		231 :
			REF <= 23'b0001101_0100011010101010;	// 1
		232 :
			REF <= 23'b0001100_0100011000100100;	// 0
		233 :
			REF <= 23'b0001100_0100011000100100;	// 1
		234 :
			REF <= 23'b0001011_0100010110011110;	// 0
		235 :
			REF <= 23'b0001011_0100010110011110;	// 1
		236 :
			REF <= 23'b0001010_0100010100011001;	// 0
		237 :
			REF <= 23'b0001010_0100010100011001;	// 1
		238 :
			REF <= 23'b0001001_0100010010010100;	// 0
		239 :
			REF <= 23'b0001001_0100010010010100;	// 1
		240 :
			REF <= 23'b0001000_0100010000010000;	// 1
		241 :
			REF <= 23'b0000111_0100001110001100;	// 0
		242 :
			REF <= 23'b0000111_0100001110001100;	// 1
		243 :
			REF <= 23'b0000110_0100001100001001;	// 0
		244 :
			REF <= 23'b0000110_0100001100001001;	// 1
		245 :
			REF <= 23'b0000101_0100001010000110;	// 0
		246 :
			REF <= 23'b0000101_0100001010000110;	// 1
		247 :
			REF <= 23'b0000100_0100001000000100;	// 0
		248 :
			REF <= 23'b0000100_0100001000000100;	// 1
		249 :
			REF <= 23'b0000011_0100000110000010;	// 0
		250 :
			REF <= 23'b0000011_0100000110000010;	// 1
		251 :
			REF <= 23'b0000010_0100000100000001;	// 0
		252 :
			REF <= 23'b0000010_0100000100000001;	// 1
		253 :
			REF <= 23'b0000001_0100000010000000;	// 0
		254 :
			REF <= 23'b0000001_0100000010000000;	// 1
		255 :
			REF <= 23'b0000000_0100000000000000;	// 256
	endcase
end

endmodule
